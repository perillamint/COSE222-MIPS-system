`include "simparams.vh"

// Hazard detection unit

module hdu(input clk, input reset);
endmodule // hdu
