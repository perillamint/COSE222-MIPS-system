parameter res_x = 320;
parameter res_y = 200;
parameter fbsize = res_x * res_y / 8;
