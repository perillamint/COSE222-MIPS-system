`timescale 1ns/1ps
`define mydelay 1
